`timescale 1ns/1ns 
import uvm_pkg::*; 
`include "uvm_macros.svh" 
//-------------------------------------------------------- 
//Include Files 
//-------------------------------------------------------- 
`include "interface.sv" 
`include "sequence_item.sv" 
`include "sequence.sv" 
`include "sequencer.sv" 
`include "driver.sv" 
`include "monitor.sv" 
`include "agent.sv" 
`include "scoreboard.sv" 
`include "environment.sv" 
`include "test.sv" 
module top; 
//-------------------------------------------------------- 
//Instantiation 
//-------------------------------------------------------- 
logic clock; 
alu_interface intf(.clock(clock)); 
alu dut( 
.clock(intf.clock), 
.reset(intf.reset), 
.A(intf.a), 
.B(intf.b), 
.ALU_Sel(intf.op_code), 
.ALU_Out(intf.result), 
.CarryOut(intf.carry_out) 
); 
                                                                                                                                                         //-------------------------------------------------------- 
  //Interface Setting 
  //-------------------------------------------------------- 
  initial begin 
    uvm_config_db #(virtual alu_interface)::set(null, "*", "vif", intf ); 
 
  end 
   
   
   
  //-------------------------------------------------------- 
  //Start The Test 
  //-------------------------------------------------------- 
  initial begin 
    run_test("alu_test"); 
  end 
   
   
  //-------------------------------------------------------- 
  //Clock Generation 
  //-------------------------------------------------------- 
  initial begin 
    clock = 0; 
    #5; 
    forever begin 
      clock = ~clock; 
      #2; 
    end 
  end 
   
   
  //-------------------------------------------------------- 
  //Maximum Simulation Time 
  //-------------------------------------------------------- 
  initial begin 
    #5000; 
    $display("Sorry! Ran out of clock cycles!"); 
    $finish(); 
  end 
   
   
  //-------------------------------------------------------- 
  //Generate Waveforms 
  //-------------------------------------------------------- 
  initial begin 
    $dumpfile("d.vcd"); 
    $dumpvars(); 
  end 
   
   
   
endmodule: top
